// L1_WEIGHTS
localparam [7:0] L1_WEIGHTS[0:7] = '{
  8'b10100000,
  8'b01000001,
  8'b01111010,
  8'b00011000,
  8'b11101101,
  8'b10110111,
  8'b01100111,
  8'b00111010
};
// L2_WEIGHTS
localparam [7:0] L2_WEIGHTS[0:3] = '{
  8'b11111001,
  8'b01100010,
  8'b11110111,
  8'b00001111
};
