// L1_WEIGHTS
localparam [7:0] L1_WEIGHTS[0:7] = '{
  8'b11010111,
  8'b10000110,
  8'b11111001,
  8'b10001111,
  8'b11100100,
  8'b10101001,
  8'b11101000,
  8'b10111000
};

// L2_WEIGHTS
localparam [7:0] L2_WEIGHTS[0:3] = '{
  8'b01010001,
  8'b00000110,
  8'b00001001,
  8'b10011010
};
